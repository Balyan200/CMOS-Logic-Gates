magic
tech scmos
timestamp 1754233407
<< nwell >>
rect -13 -19 15 14
<< ntransistor >>
rect 0 -42 2 -37
<< ptransistor >>
rect 0 -13 2 0
<< ndiffusion >>
rect -2 -42 0 -37
rect 2 -42 4 -37
<< pdiffusion >>
rect -2 -4 0 0
rect -6 -7 0 -4
rect -2 -11 0 -7
rect -6 -13 0 -11
rect 2 -4 4 0
rect 2 -7 8 -4
rect 2 -11 4 -7
rect 2 -13 8 -11
<< ndcontact >>
rect -6 -42 -2 -37
rect 4 -42 8 -37
<< pdcontact >>
rect -6 -4 -2 0
rect -6 -11 -2 -7
rect 4 -4 8 0
rect 4 -11 8 -7
<< psubstratepcontact >>
rect -13 -50 -9 -46
rect 4 -50 8 -46
<< nsubstratencontact >>
rect -8 7 -4 11
rect 4 7 8 11
<< polysilicon >>
rect 0 0 2 4
rect 0 -24 2 -13
rect -4 -25 2 -24
rect 0 -34 2 -30
rect -4 -35 2 -34
rect 0 -37 2 -35
rect 0 -45 2 -42
<< polycontact >>
rect -4 -24 0 -20
rect -4 -34 0 -30
<< metal1 >>
rect -13 11 15 12
rect -13 7 -8 11
rect -4 7 4 11
rect 8 7 15 11
rect -13 6 15 7
rect -6 0 -1 6
rect -2 -4 -1 0
rect -6 -7 -1 -4
rect -2 -11 -1 -7
rect -6 -13 -1 -11
rect 3 -4 4 0
rect 3 -7 8 -4
rect 3 -11 4 -7
rect -4 -25 0 -24
rect -15 -29 0 -25
rect -4 -30 0 -29
rect 3 -25 8 -11
rect 3 -29 17 -25
rect 3 -37 8 -29
rect -2 -42 -1 -37
rect 3 -42 4 -37
rect -6 -46 -1 -42
rect -16 -50 -13 -46
rect -9 -50 4 -46
rect 8 -50 17 -46
<< labels >>
rlabel metal1 -13 -27 -13 -27 3 in
rlabel psubstratepcontact -12 -48 -12 -48 2 gnd
rlabel metal1 13 -27 13 -27 7 out
rlabel metal1 -1 9 -1 9 5 vdd
<< end >>
